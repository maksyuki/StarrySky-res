`timescale 1ns / 1ps

`define chiplink_data_w 8

module chiplink_ctrl (
    input                             clk,
    input                             resetn,
    output                            chiplink_rx_clk,
    output                            chiplink_rx_rst,
    output                            chiplink_rx_send,
    output [`chiplink_data_w - 1 : 0] chiplink_rx_data,

    input                             chiplink_tx_clk,
    input                             chiplink_tx_rst,
    input                             chiplink_tx_send,
    input  [`chiplink_data_w - 1 : 0] chiplink_tx_data,
    output                            chiplink_cpu_int,

    input         io_axi4_0_awready,
    output        io_axi4_0_awvalid,
    output [ 3:0] io_axi4_0_awid,
    output [31:0] io_axi4_0_awaddr,
    output [ 7:0] io_axi4_0_awlen,
    output [ 2:0] io_axi4_0_awsize,
    output [ 1:0] io_axi4_0_awburst,
    input         io_axi4_0_wready,
    output        io_axi4_0_wvalid,
    output [63:0] io_axi4_0_wdata,
    output [ 7:0] io_axi4_0_wstrb,
    output        io_axi4_0_wlast,
    output        io_axi4_0_bready,
    input         io_axi4_0_bvalid,
    input  [ 3:0] io_axi4_0_bid,
    input  [ 1:0] io_axi4_0_bresp,
    input         io_axi4_0_arready,
    output        io_axi4_0_arvalid,
    output [ 3:0] io_axi4_0_arid,
    output [31:0] io_axi4_0_araddr,
    output [ 7:0] io_axi4_0_arlen,
    output [ 2:0] io_axi4_0_arsize,
    output [ 1:0] io_axi4_0_arburst,
    output        io_axi4_0_rready,
    input         io_axi4_0_rvalid,
    input  [ 3:0] io_axi4_0_rid,
    input  [63:0] io_axi4_0_rdata,
    input  [ 1:0] io_axi4_0_rresp,
    input         io_axi4_0_rlast
);

  wire [31:0] aw_addr;
  wire [31:0] ar_addr;
  //chiplink sim connect to dual chiplink
  FPGA_ChiplinkBridge u_FPGA_ChiplinkBridge (
      .clock                         (clk),
      .reset                         (~resetn),
      .fpga_io_c2b_clk               (chiplink_rx_clk),
      .fpga_io_c2b_rst               (chiplink_rx_rst),
      .fpga_io_c2b_send              (chiplink_rx_send),
      .fpga_io_c2b_data              (chiplink_rx_data),
      .fpga_io_b2c_clk               (chiplink_tx_clk),
      .fpga_io_b2c_rst               (chiplink_tx_rst),
      .fpga_io_b2c_send              (chiplink_tx_send),
      .fpga_io_b2c_data              (chiplink_tx_data),
      //mem
      .mem_axi4_0_awready            (io_axi4_0_awready),
      .mem_axi4_0_awvalid            (io_axi4_0_awvalid),
      .mem_axi4_0_awid               (io_axi4_0_awid),
      .mem_axi4_0_awaddr             (aw_addr),
      .mem_axi4_0_awlen              (io_axi4_0_awlen),
      .mem_axi4_0_awsize             (io_axi4_0_awsize),
      .mem_axi4_0_awburst            (io_axi4_0_awburst),
      .mem_axi4_0_wready             (io_axi4_0_wready),
      .mem_axi4_0_wvalid             (io_axi4_0_wvalid),
      .mem_axi4_0_wdata              (io_axi4_0_wdata),
      .mem_axi4_0_wstrb              (io_axi4_0_wstrb),
      .mem_axi4_0_wlast              (io_axi4_0_wlast),
      .mem_axi4_0_bready             (io_axi4_0_bready),
      .mem_axi4_0_bvalid             (io_axi4_0_bvalid),
      .mem_axi4_0_bid                (io_axi4_0_bid),
      .mem_axi4_0_bresp              (io_axi4_0_bresp),
      .mem_axi4_0_arready            (io_axi4_0_arready),
      .mem_axi4_0_arvalid            (io_axi4_0_arvalid),
      .mem_axi4_0_arid               (io_axi4_0_arid),
      .mem_axi4_0_araddr             (ar_addr),
      .mem_axi4_0_arlen              (io_axi4_0_arlen),
      .mem_axi4_0_arsize             (io_axi4_0_arsize),
      .mem_axi4_0_arburst            (io_axi4_0_arburst),
      .mem_axi4_0_rready             (io_axi4_0_rready),
      .mem_axi4_0_rvalid             (io_axi4_0_rvalid),
      .mem_axi4_0_rid                (io_axi4_0_rid),
      .mem_axi4_0_rdata              (io_axi4_0_rdata),
      .mem_axi4_0_rresp              (io_axi4_0_rresp),
      .mem_axi4_0_rlast              (io_axi4_0_rlast),
      //dma
      .slave_axi4_mem_0_awready(),
      .slave_axi4_mem_0_awvalid(1'b0),
      .slave_axi4_mem_0_awid(4'b0),
      .slave_axi4_mem_0_awaddr(32'b0),
      .slave_axi4_mem_0_awlen(8'b0),
      .slave_axi4_mem_0_awsize(3'b0),
      .slave_axi4_mem_0_awburst(2'b0),
      .slave_axi4_mem_0_wready(),
      .slave_axi4_mem_0_wvalid(1'b0),
      .slave_axi4_mem_0_wdata(64'b0),
      .slave_axi4_mem_0_wstrb(8'b0),
      .slave_axi4_mem_0_wlast(1'b0),
      .slave_axi4_mem_0_bready(1'b0),
      .slave_axi4_mem_0_bvalid(),
      .slave_axi4_mem_0_bid(),
      .slave_axi4_mem_0_bresp(),
      .slave_axi4_mem_0_arready(),
      .slave_axi4_mem_0_arvalid(1'b0),
      .slave_axi4_mem_0_arid(4'b0),
      .slave_axi4_mem_0_araddr(32'b0),
      .slave_axi4_mem_0_arlen(8'b0),
      .slave_axi4_mem_0_arsize(3'b0),
      .slave_axi4_mem_0_arburst(2'b0),
      .slave_axi4_mem_0_rready(1'b0),
      .slave_axi4_mem_0_rvalid(),
      .slave_axi4_mem_0_rid(),
      .slave_axi4_mem_0_rdata(),
      .slave_axi4_mem_0_rresp(),
      .slave_axi4_mem_0_rlast()
  );
  
  assign io_axi4_0_awaddr = aw_addr - 32'h8000_0000 + 32'h10_0000;
  assign io_axi4_0_araddr = ar_addr - 32'h8000_0000 + 32'h10_0000;
  assign chiplink_cpu_int = 1'b0;
endmodule
